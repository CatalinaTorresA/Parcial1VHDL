library verilog;
use verilog.vl_types.all;
entity CONPAR_vlg_vec_tst is
end CONPAR_vlg_vec_tst;
